library verilog;
use verilog.vl_types.all;
entity load_vlg_vec_tst is
end load_vlg_vec_tst;
