library verilog;
use verilog.vl_types.all;
entity load_vlg_check_tst is
    port(
        pulse_out       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end load_vlg_check_tst;
